module reference_search_area_centre(input [5:0] counter, output [6:0] x_centre_reference, y_centre_reference);
wire [6:0] x_centre[0:35];
wire [6:0] y_centre[0:35];
assign x_centre[0]=16;
assign x_centre[1]=16;
assign x_centre[2]=16;
assign x_centre[3]=16;
assign x_centre[4]=16;
assign x_centre[5]=16;
assign x_centre[6]=24;
assign x_centre[7]=24;
assign x_centre[8]=24;
assign x_centre[9]=24;
assign x_centre[10]=24;
assign x_centre[11]=24;
assign x_centre[12]=40;
assign x_centre[13]=40;
assign x_centre[14]=40;
assign x_centre[15]=40;
assign x_centre[16]=40;
assign x_centre[17]=40;
assign x_centre[18]=56;
assign x_centre[19]=56;
assign x_centre[20]=56;
assign x_centre[21]=56;
assign x_centre[22]=56;
assign x_centre[23]=56;
assign x_centre[24]=72;
assign x_centre[25]=72;
assign x_centre[26]=72;
assign x_centre[27]=72;
assign x_centre[28]=72;
assign x_centre[29]=72;
assign x_centre[30]=80;
assign x_centre[31]=80;
assign x_centre[32]=80;
assign x_centre[33]=80;
assign x_centre[34]=80;
assign x_centre[35]=80;

assign y_centre[0]=16;
assign y_centre[1]=24;
assign y_centre[2]=40;
assign y_centre[3]=56;
assign y_centre[4]=72;
assign y_centre[5]=80;
assign y_centre[6]=16;
assign y_centre[7]=24;
assign y_centre[8]=40;
assign y_centre[9]=56;
assign y_centre[10]=72;
assign y_centre[11]=80;
assign y_centre[12]=16;
assign y_centre[13]=24;
assign y_centre[14]=40;
assign y_centre[15]=56;
assign y_centre[16]=72;
assign y_centre[17]=80;
assign y_centre[18]=16;
assign y_centre[19]=24;
assign y_centre[20]=40;
assign y_centre[21]=56;
assign y_centre[22]=72;
assign y_centre[23]=80;
assign y_centre[24]=16;
assign y_centre[25]=24;
assign y_centre[26]=40;
assign y_centre[27]=56;
assign y_centre[28]=72;
assign y_centre[29]=80;
assign y_centre[30]=16;
assign y_centre[31]=24;
assign y_centre[32]=40;
assign y_centre[33]=56;
assign y_centre[34]=72;
assign y_centre[35]=80;

//fetching the centre coordinates from the register file
assign x_centre_reference=x_centre[counter];
assign y_centre_reference=y_centre[counter];

endmodule
